module ICache();

endmodule
