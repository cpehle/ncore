module CSRFile(input clk);

endmodule
