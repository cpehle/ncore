module RRArbiter();

endmodule
