`include "Bundle.sv"
module Alu(
           input Bundle::AluIn alu_in,
           output Bundle::AluOut alu_out
);


endmodule; // Alu
