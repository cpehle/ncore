module DutReplayBuffer();

endmodule // DutReplayBuffer
// Local Variables:
// verilog-library-directories:("." "../src/")
// End:
