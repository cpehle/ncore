module BranchTargetBuffer(
			  BTBRequest req,			
);
endmodule // BranchTargetBuffer

module BranchHistoryTable();
endmodule // BranchHistoryTable

