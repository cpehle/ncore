module BranchHistoryTable();
endmodule
