///@file RouterOutput.sv
///@author Christian Pehle
///@brief
module RouterOutput();

endmodule
