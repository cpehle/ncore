module WriteBack();


endmodule
