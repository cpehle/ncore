module Memory();


endmodule
