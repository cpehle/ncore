module InstructionFetchUnit();

   genvar i;
   generate
      


   endgenerate

endmodule
