module test_axi_register(input clk);

   

   
endmodule
