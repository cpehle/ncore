module RRArbiter #(parameter int width = 2) ();

endmodule
