// file: TLB
//
// Translation Lookaside Buffer
module TLB();
endmodule
