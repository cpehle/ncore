`include "Bundle.sv"
module BranchTargetBuffer(
			  input Bundle::BTBRequest req
);

endmodule // BranchTargetBuffer


