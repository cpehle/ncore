module RegisterFile();
endmodule; // RegisterFile
