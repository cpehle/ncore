`ifndef _Instructions
`define _Instructions
package Instructions;
`define MCRF       32'b100110???????????????0000000000?
`define BCLR       32'b100110???????????????1000000000?
`define CRNOR      32'b100110???????????????1000010000?
`define RFMCI      32'b100110???????????????1001100000?
`define RFI        32'b100110???????????????1100100000?
`define RFCI       32'b100110???????????????1100110000?
`define CRXOR      32'b100110???????????????1100000100?
`define CRNAND     32'b100110???????????????1110000100?
`define CRANDC     32'b100110???????????????1000000100?
`define CREQV      32'b100110???????????????1001000010?
`define CRAND      32'b100110???????????????1000000010?
`define CRORC      32'b100110???????????????1101000010?
`define CROR       32'b100110???????????????1110000010?
`define BCCTR      32'b100110???????????????1000010000?
`define SUBFC      32'b111110????????????????100000000?
`define ADDC       32'b111110????????????????101000000?
`define MULHWU     32'b111110????????????????101100000?
`define SUBF       32'b111110????????????????101000000?
`define MULHW      32'b111110????????????????100101100?
`define NEG        32'b111110????????????????110100000?
`define SUBFE      32'b111110????????????????100010000?
`define ADDE       32'b111110????????????????100010100?
`define SUBFZE     32'b111110????????????????110010000?
`define ADDZE      32'b111110????????????????110010100?
`define SUBFME     32'b111110????????????????111010000?
`define ADDME      32'b111110????????????????111010100?
`define MULLW      32'b111110????????????????111010110?
`define ADD        32'b111110????????????????100001010?
`define DIVWU      32'b111110????????????????111001011?
`define DIVW       32'b111110????????????????111101011?
`define CMP        32'b111110???????????????0000000000?
`define TW         32'b111110???????????????1000000000?
`define LWZX       32'b111110???????????????1011100000?
`define SLW        32'b111110???????????????1100000000?
`define CNTLZW     32'b111110???????????????1101000000?
`define AND        32'b111110???????????????1110000000?
`define CMPL       32'b111110???????????????1000000000?
`define NVEM       32'b111110???????????????1100000000?
`define NVES       32'b111110???????????????1100010000?
`define NVEMTL     32'b111110???????????????1100100000?
`define LWZUX      32'b111110???????????????1101110000?
`define ANDC       32'b111110???????????????1111000000?
`define WAIT       32'b111110???????????????1111100000?
`define MFMSR      32'b111110???????????????1010011000?
`define LBZX       32'b111110???????????????1010111000?
`define LBZUX      32'b111110???????????????1110111000?
`define POPCB      32'b111110???????????????1111010000?
`define NOR        32'b111110???????????????1111100000?
`define MTMSR      32'b111110???????????????1001001000?
`define STWX       32'b111110???????????????1001011100?
`define PRTYW      32'b111110???????????????1001101000?
`define STWUX      32'b111110???????????????1011011100?
`define STBX       32'b111110???????????????1101011100?
`define STBUX      32'b111110???????????????1111011100?
`define LHZX       32'b111110???????????????1000101110?
`define EQV        32'b111110???????????????1000111000?
`define ECIWX      32'b111110???????????????1001101100?
`define LHZUX      32'b111110???????????????1001101110?
`define XOR        32'b111110???????????????1001111000?
`define POPCW      32'b111110???????????????1011110100?
`define LHAX       32'b111110???????????????1010101110?
`define LHAUX      32'b111110???????????????1011101110?
`define STHX       32'b111110???????????????1100101110?
`define ORC        32'b111110???????????????1100111000?
`define ECOWX      32'b111110???????????????1101101100?
`define STHUX      32'b111110???????????????1101101110?
`define OR         32'b111110???????????????1101111000?
`define NAND       32'b111110???????????????1110111000?
`define SRW        32'b111110???????????????1000011000?
`define TWI        32'b110000??????????????????????????
`define MULLI      32'b111000??????????????????????????
`define SUBFIC     32'b100000??????????????????????????
`define CMPLI      32'b101000??????????????????????????
`define CMPI       32'b101100??????????????????????????
`define ADDIC      32'b110000??????????????????????????
`define ADDI       32'b111000??????????????????????????
`define ADDIS      32'b111100??????????????????????????
`define BC         32'b100000??????????????????????????
`define BRANCH     32'b100100??????????????????????????
`define RLWIMI     32'b101000??????????????????????????
`define RLWINM     32'b101010??????????????????????????
`define RLWNM      32'b101110??????????????????????????
`define ORI        32'b110000??????????????????????????
`define ORIS       32'b110010??????????????????????????
`define XORI       32'b110100??????????????????????????
`define XORIS      32'b110110??????????????????????????
`define ANDI       32'b111000??????????????????????????
`define ANDIS      32'b111010??????????????????????????
`define LWZ        32'b100000??????????????????????????
`define LWZU       32'b100001??????????????????????????
`define LBZ        32'b100010??????????????????????????
`define LBZU       32'b100011??????????????????????????
`define STW        32'b100100??????????????????????????
`define STWU       32'b100101??????????????????????????
`define STB        32'b100110??????????????????????????
`define STBU       32'b100111??????????????????????????
`define LHZ        32'b101000??????????????????????????
`define LHZU       32'b101001??????????????????????????
`define LHA        32'b101010??????????????????????????
`define LHAU       32'b101011??????????????????????????
`define STH        32'b101100??????????????????????????
`define STHU       32'b101101??????????????????????????
`define LMW        32'b101110??????????????????????????
`define STMW       32'b101111??????????????????????????
endpackage
`endif
