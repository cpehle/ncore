`ifndef _Instructions
`define _Instructions
package Instructions;
`define MCRF       32'b10011????????????????0??????????
`define BCLR       32'b10011????????????????10000??????
`define CRNOR      32'b10011????????????????100001?????
`define RFMCI      32'b10011????????????????100110?????
`define RFI        32'b10011????????????????110010?????
`define RFCI       32'b10011????????????????110011?????
`define CRXOR      32'b10011????????????????11000001???
`define CRNAND     32'b10011????????????????11100001???
`define CRANDC     32'b10011????????????????10000001???
`define CREQV      32'b10011????????????????100100001??
`define CRAND      32'b10011????????????????100000001??
`define CRORC      32'b10011????????????????110100001??
`define CROR       32'b10011????????????????111000001??
`define BCCTR      32'b10011????????????????1000010000?
`define SUBFC      32'b11111?????????????????1000??????
`define ADDC       32'b11111?????????????????1010??????
`define MULHWU     32'b11111?????????????????1011??????
`define SUBF       32'b11111?????????????????101000????
`define MULHW      32'b11111?????????????????1001011???
`define NEG        32'b11111?????????????????1101000???
`define SUBFE      32'b11111?????????????????10001000??
`define ADDE       32'b11111?????????????????10001010??
`define SUBFZE     32'b11111?????????????????11001000??
`define ADDZE      32'b11111?????????????????11001010??
`define SUBFME     32'b11111?????????????????11101000??
`define ADDME      32'b11111?????????????????11101010??
`define MULLW      32'b11111?????????????????11101011??
`define ADD        32'b11111?????????????????100001010?
`define DIVWU      32'b11111?????????????????111001011?
`define DIVW       32'b11111?????????????????111101011?
`define CMP        32'b11111????????????????0??????????
`define TW         32'b11111????????????????100????????
`define LWZX       32'b11111????????????????10111??????
`define SLW        32'b11111????????????????11000??????
`define CNTLZW     32'b11111????????????????11010??????
`define AND        32'b11111????????????????11100??????
`define CMPL       32'b11111????????????????100000?????
`define NVEM       32'b11111????????????????110000?????
`define NVES       32'b11111????????????????110001?????
`define NVEMTL     32'b11111????????????????110010?????
`define LWZUX      32'b11111????????????????110111?????
`define ANDC       32'b11111????????????????111100?????
`define WAIT       32'b11111????????????????111110?????
`define MFMSR      32'b11111????????????????1010011????
`define LBZX       32'b11111????????????????1010111????
`define LBZUX      32'b11111????????????????1110111????
`define POPCB      32'b11111????????????????1111010????
`define NOR        32'b11111????????????????1111100????
`define MTMSR      32'b11111????????????????10010010???
`define STWX       32'b11111????????????????10010111???
`define PRTYW      32'b11111????????????????10011010???
`define STWUX      32'b11111????????????????10110111???
`define STBX       32'b11111????????????????11010111???
`define STBUX      32'b11111????????????????11110111???
`define LHZX       32'b11111????????????????100010111??
`define EQV        32'b11111????????????????100011100??
`define ECIWX      32'b11111????????????????100110110??
`define LHZUX      32'b11111????????????????100110111??
`define XOR        32'b11111????????????????100111100??
`define POPCW      32'b11111????????????????101111010??
`define LHAX       32'b11111????????????????101010111??
`define LHAUX      32'b11111????????????????101110111??
`define STHX       32'b11111????????????????110010111??
`define ORC        32'b11111????????????????110011100??
`define ECOWX      32'b11111????????????????110110110??
`define STHUX      32'b11111????????????????110110111??
`define OR         32'b11111????????????????110111100??
`define NAND       32'b11111????????????????111011100??
`define SRW        32'b11111????????????????1000011000?
`define TWI        32'b11??????????????????????????????
`define MULLI      32'b111?????????????????????????????
`define SUBFIC     32'b1000????????????????????????????
`define CMPLI      32'b1010????????????????????????????
`define CMPI       32'b1011????????????????????????????
`define ADDIC      32'b1100????????????????????????????
`define ADDI       32'b1110????????????????????????????
`define ADDIS      32'b1111????????????????????????????
`define BC         32'b10000???????????????????????????
`define BRANCH     32'b10010???????????????????????????
`define RLWIMI     32'b10100???????????????????????????
`define RLWINM     32'b10101???????????????????????????
`define RLWNM      32'b10111???????????????????????????
`define ORI        32'b11000???????????????????????????
`define ORIS       32'b11001???????????????????????????
`define XORI       32'b11010???????????????????????????
`define XORIS      32'b11011???????????????????????????
`define ANDI       32'b11100???????????????????????????
`define ANDIS      32'b11101???????????????????????????
`define LWZ        32'b100000??????????????????????????
`define LWZU       32'b100001??????????????????????????
`define LBZ        32'b100010??????????????????????????
`define LBZU       32'b100011??????????????????????????
`define STW        32'b100100??????????????????????????
`define STWU       32'b100101??????????????????????????
`define STB        32'b100110??????????????????????????
`define STBU       32'b100111??????????????????????????
`define LHZ        32'b101000??????????????????????????
`define LHZU       32'b101001??????????????????????????
`define LHA        32'b101010??????????????????????????
`define LHAU       32'b101011??????????????????????????
`define STH        32'b101100??????????????????????????
`define STHU       32'b101101??????????????????????????
`define LMW        32'b101110??????????????????????????
`define STMW       32'b101111??????????????????????????
endpackage
`endif
