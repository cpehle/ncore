`ifndef _Instructions
`define _Instructions
package Instructions;
`define BEQ 32'b?????????????????000?????1100011
`define BNE 32'b?????????????????001?????1100011
`define BLT 32'b?????????????????100?????1100011
`define BGE 32'b?????????????????101?????1100011
`define BLTU 32'b?????????????????110?????1100011
`define BGEU 32'b?????????????????111?????1100011
`define JALR 32'b?????????????????000?????1100111
`define JAL 32'b?????????????????????????1101111
`define LUI 32'b?????????????????????????0110111
`define AUIPC 32'b?????????????????????????0010111
`define ADDI 32'b?????????????????000?????0010011
`define SLLI 32'b000000???????????001?????0010011
`define SLTI 32'b?????????????????010?????0010011
`define SLTIU 32'b?????????????????011?????0010011
`define XORI 32'b?????????????????100?????0010011
`define SRLI 32'b000000???????????101?????0010011
`define SRAI 32'b010000???????????101?????0010011
`define ORI 32'b?????????????????110?????0010011
`define ANDI 32'b?????????????????111?????0010011
`define ADD 32'b0000000??????????000?????0110011
`define SUB 32'b0100000??????????000?????0110011
`define SLL 32'b0000000??????????001?????0110011
`define SLT 32'b0000000??????????010?????0110011
`define SLTU 32'b0000000??????????011?????0110011
`define XOR 32'b0000000??????????100?????0110011
`define SRL 32'b0000000??????????101?????0110011
`define SRA 32'b0100000??????????101?????0110011
`define OR 32'b0000000??????????110?????0110011
`define AND 32'b0000000??????????111?????0110011
`define ADDIW 32'b?????????????????000?????0011011
`define SLLIW 32'b0000000??????????001?????0011011
`define SRLIW 32'b0000000??????????101?????0011011
`define SRAIW 32'b0100000??????????101?????0011011
`define ADDW 32'b0000000??????????000?????0111011
`define SUBW 32'b0100000??????????000?????0111011
`define SLLW 32'b0000000??????????001?????0111011
`define SRLW 32'b0000000??????????101?????0111011
`define SRAW 32'b0100000??????????101?????0111011
`define LB 32'b?????????????????000?????0000011
`define LH 32'b?????????????????001?????0000011
`define LW 32'b?????????????????010?????0000011
`define LD 32'b?????????????????011?????0000011
`define LBU 32'b?????????????????100?????0000011
`define LHU 32'b?????????????????101?????0000011
`define LWU 32'b?????????????????110?????0000011
`define SB 32'b?????????????????000?????0100011
`define SH 32'b?????????????????001?????0100011
`define SW 32'b?????????????????010?????0100011
`define SD 32'b?????????????????011?????0100011
`define FENCE 32'b?????????????????000?????0001111
`define FENCE_I 32'b?????????????????001?????0001111

`define SCALL 32'b00000000000000000000000001110011
`define SBREAK 32'b00000000000100000000000001110011
`define SRET 32'b00010000000000000000000001110011
`define WFI 32'b00010000001000000000000001110011

`define MRTS 32'b00110000010100000000000001110011

`define CSRRW 32'b?????????????????001?????1110011
`define CSRRS 32'b?????????????????010?????1110011
`define CSRRC 32'b?????????????????011?????1110011
`define CSRRWI 32'b?????????????????101?????1110011
`define CSRRSI 32'b?????????????????110?????1110011
`define CSRRCI 32'b?????????????????111?????1110011
endpackage
`endif
