module TraceCache(
);
endmodule // TraceCache
