package DMA;

endpackage
