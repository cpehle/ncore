module InstructionFetch();

endmodule
