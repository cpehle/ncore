module Alu();
endmodule; // Alu
