module BreakpointUnit(input clk);
endmodule
