

module DutInstructionDecode();


endmodule
