module TraceCache();
endmodule
